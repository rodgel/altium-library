.SUBCKT GT20D101 71 72 74
*     TERMINALS:  C  G  E
*  250 Volt  20 Amp  17.2NS  N-Channel IGBT  09-15-1992
Q1  83 81 85     QOUT
M1  81 82 83 83  MFIN L=1U W=1U
DSD 83 81  DO
DBE 85 81  DE
RC  85 71  66.5M
RE  83 73  6.65M
RG  72 82  23.2
CGE 82 83  1.33N
CGC 82 71  1P
EGD 91  0 82 81  1
VFB 93  0  0
FFB 82 81  VFB  1
CGD 92 93  457P
R1  92  0  1
D1  91 92  DLIM
DHV 94 93  DR
R2  91 94  1
D2  94  0  DLIM
LE  73 74  7.5N
.MODEL QOUT PNP (IS=10.1F NF=1.2 BF=5.1 CJE=2.25N TF=17.2N XTB=1.3)
.MODEL MFIN NMOS (LEVEL=3 VMAX=221K THETA=80M ETA=4.81M VTO=3 KP=1.29)
.MODEL DR D (IS=1.01F CJO=457P VJ=1 M=.82)
.MODEL DO D (IS=1.01F BV=250 CJO=1.79N VJ=1 M=.7)
.MODEL DE D (IS=1.01F BV=14.3 N=2)
.MODEL DLIM D (IS=100N)
.ENDS 